`ifndef CONSTANTS
`define CONSTANTS

`define OPCODE_I 7'b0010011
`define OPCODE_R 7'b1100011

`define FUNC3_ADD 3'b000
`define FUNC3_OR 3'b110
`define FUNC3_AND 3'b111

`define ALU_ADD	3'b000
`define ALU_OR		3'b001
`define ALU_AND	3'b010

`endif