`ifndef CONSTANTS
`define CONSTANTS

`define FUNC3_ADD 5'b000
`define F_SUB 5'b00010

`endif