`ifndef CONSTANTS
`define CONSTANTS

`define F_ADD 5'b00001
`define F_SUB 5'b00010

`endif